library verilog;
use verilog.vl_types.all;
entity ClockTop_tb is
end ClockTop_tb;
